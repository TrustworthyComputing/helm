module adder(G11, G12, G14);
  wire 00, 01, 02, 03, 04, 05, 06, 07, 08, 09, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 56, 57, 58;
  input [7:0] G11;
  input [7:0] G12;
  output [7:0] G14;
  lut lut_gate1(0x8778, G12[1], G11[1], G12[0], G11[0], G14[1]);
  lut lut_gate2(0xf880077f077ff880, G12[2], G11[2], G12[1], G11[1], G12[0], G11[0], G14[2]);
  lut lut_gate3(0x0317173f173f173f, G11[0], G12[0], G12[1], G12[2], G11[2], G11[1], 56);
  lut lut_gate4(0x69, G12[3], G11[3], 56, G14[3]);
  lut lut_gate5(3559599060, G12[4], G11[4], G12[3], G11[3], 56, G14[4]);
  lut lut_gate6(53160767, G12[3], G11[3], G12[4], G11[4], 56, 57);
  lut lut_gate7(0x69, G12[5], G11[5], 57, G14[5]);
  lut lut_gate8(3559599060, G12[6], G11[6], G12[5], G11[5], 57, G14[6]);
  lut lut_gate9(0x6, G12[7], G11[7], 58);
  lut lut_gate10(0x032b2b3ffc, 58, G12[5], G11[5], G12[6], G11[6], 57, G14[7]);
  lut lut_gate11(0x6, G12[0], G11[0], G14[0]);

endmodule
